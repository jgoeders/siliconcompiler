(* blackbox *)
module bit_or (
  input clk,
  input nrst,

  input a,
  input b,

  output reg y
);
endmodule
