(* blackbox *)
module bit_and (
  input clk,
  input nrst,

  input a,
  input b,

  output reg y
);
endmodule
